


package SPI_pkg;


 import uvm_pkg::*;
 
 `include "uvm_macros.svh"
  

  `include "SPI_seq_item.sv"
  `include "Sequence.sv"
  `include "Sequencer.sv"   
  `include "Driver.sv"  
  `include "Monitor.sv"
  `include "Coverage_collector.sv"
  `include "Agent.sv"  
  `include "Environment.sv"  
  `include "SPI_Test.sv"

 

endpackage 